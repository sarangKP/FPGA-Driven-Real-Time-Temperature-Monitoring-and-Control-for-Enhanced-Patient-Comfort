//This is a testbench and was written for testing only
module DHT11_tb(); 
	reg clk_tb; 
	wire w1_tb; 
	wire done_tb;
	wire [7:0] temp_tb;
	wire [7:0] hum_tb;
	
	reg w1r; 
	reg w1_en; 
	
	DHT11 DHT11_tb(clk_tb, w1_tb, done_tb, temp_tb, hum_tb); 
	initial begin 
			clk_tb <= 1'b0; 
			w1r <= 1'b0; 
			w1_en <= 1'b0; 
	end 
	
	always begin 
		#10
			clk_tb <= ~clk_tb; 
	end
	
	always begin 
		#21000000
			w1r <= 1'b0; 
			w1_en <= 1'b1; 
		#80000
			w1r <= 1'b1;
		#80000
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 1 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 2 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 3 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 4 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 5 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 6 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 7 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 8 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 9 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 10 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 11 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 12 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 13 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 14 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 15 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 16 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 17 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 18 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 19 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 20 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 21 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 22 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 23 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 24 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 25 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 26 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 27 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 28 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 29 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 30 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 31 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 32 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 33 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 34 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 35 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 36 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 37 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 38 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 39 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 40 = 1
			w1_en <= 1'b0; 
		#42000000
			w1r <= 1'b0; 
			w1_en <= 1'b1; 
		#80000
			w1r <= 1'b1;
		#80000
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 1 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 2 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 3 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 4 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 5 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 6 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 7 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 8 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 9 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 10 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 11 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 12 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 13 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 14 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 15 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 16 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 17 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 18 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 19 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 20 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 21 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 22 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 23 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 24 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 25 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 26 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 27 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 28 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 29 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 30 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 31 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 32 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 33 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 34 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 35 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 36 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 37 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 38 = 1
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#28000 //Data 39 = 0
			w1r <= 1'b0;	
		#50000 
			w1r <= 1'b1;		
		#70000 //Data 40 = 1
			w1_en <= 1'b0;
		#21000000
			w1_en <= 1'b0;
	end 
	
	assign w1_tb = w1_en ? w1r : 1'bZ;  
	
endmodule 

